
module pc(input [63:0]loc,output [63:0]Loc);

assign Loc=loc;

endmodule

